module example_coverage(
    input clk,
    input reset_n
);
endmodule: example_coverage