module example(
    input clk,
    input reset_n
);
endmodule: example